* main circuit file
.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 1

* MUX test
Vdd Vdd 0 supplyVoltage

Va A 0 0
Vb B 0 0
Vc C 0 supplyVoltage

V_D D 0 PULSE(0, supplyVoltage, 13n, 1n, 1n, 7n, 20n)
V_CLK CLK 0 PULSE(0, supplyVoltage, 0n, 1n, 1n, 10n, 20n)

xD_LATCH D NOT_Q CLK Vdd 0 D_LATCH
xNOT NOT_Q Q Vdd 0 NOT


* plots
.plot v(Q) v(D) v(CLK)
.plot v(Q)
.plot v(CLK)
.plot v(D)

* analasys
.tran 1n 60n
module inverter(
    input a,
    output y
);

not(y,a);

endmodule
[aimspice]
[description]
422
* main circuit file
*.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 1

* circuit
Vdd Vdd 0 supplyVoltage

R1 OUT 0 1k

V_CONTROL CONTROL 0 PULSE(0, 0, 0, 2n, 2n, 50n, 60n)
V_IN IN 0 PULSE(0, supplyVoltage, 10n, 2n, 2n, 10n, 20n)

xTRANSMISSIONGATE IN OUT CONTROL Vdd 0 TRANSMISSIONGATE

* plots
.plot V(IN) V(OUT) V(CONTROL)  

* analasys
*.tran 1n 60n




[options]
1
Gmin 1e-39
[tran]
1n
60n
X
X
0
[ana]
4 0
[end]

`include "1_bit_register.v"

module eight_bit_register (output [7:0] out,input [7:0] in, input enable, input reset, input clk);

    // 8-bit register...
    
endmodule
.param L = 150n 
.param W = 150n

* NOT gate
.subckt NOT A Q Vdd Vss
   * PMOS section 
   xMP1 Q A Vdd Vdd pmos1v l=L w=W

   * NMOS section
   xMN2 Q A Vss Vss nmos1v l=L w=W
.ends NOT

* NAND gate
.subckt NAND A B Q Vdd Vss
   * PMOS section
   xMP1 Vdd A Q Vdd pmos1v l=L w=W
   xMP2 Vdd B Q Vdd pmos1v l=L w=W

   * NMOS section
   xMN1 Q B 1 1 nmos1v l=L w=W
   xMN2 1 A Vss Vss nmos1v l=L w=W
.ends NAND

* AND gate
.subckt AND A B Q Vdd Vss
   xNAND A B intermediate Vdd Vss NAND
   xNOT intermediate Q Vdd Vss NOT
.ends AND

* NOR gate 
.subckt NOR A B Q Vdd Vss
   * PMOS section
   xMP1 Vdd A 1 Vdd pmos1v l=L w=W
   xMP2 1 B Q 1 pmos1v l=L w=W

   * NMOS section
   xMN1 Q A Vss Vss nmos1v l=L w=W
   xMN2 Q B Vss Vss nmos1v l=L w=W
.ends NOR

* OR gate
.subckt OR A B Q Vdd Vss
   xNOR A B intermediate Vdd Vss NOR
   xNOT intermediate Q Vdd Vss NOT
.ends OR

* 3AND gate
.subckt 3AND A B C Q Vdd Vss
   xAND1 A B intermediate Vdd Vss AND
   xAND2 intermediate C Q Vdd Vss AND
.ends

* 3OR gate
.subckt 3OR A B C Q Vdd Vss
   xOR1 A B intermediate Vdd Vss OR
   xOR2 intermediate C Q Vdd Vss OR
.ends

* Transmission gate
.subckt TRANSMISSION_GATE IN OUT A NOT_A Vdd Vss
   * PMOS section
   xMP1 IN NOT_A OUT Vdd pmos1v l=L w=W

   * NMOS section
   xMN1 OUT A IN Vss nmos1v l=L w=W
.ends TRANSMISSION_GATE
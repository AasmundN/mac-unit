* main circuit file
.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 1

* circuit
Vdd Vdd 0 supplyVoltage

Va A 0 PULSE(0, supplyVoltage, 10n, 1n, 1n, 10n, 30n)
Vb B 0 PULSE(0, supplyVoltage, 5n, 1n, 1n, 10n, 30n)
Vc C 0 PULSE(0, supplyVoltage, 0n, 1n, 1n, 10n, 30n)

x3AND A B C Q Vdd 0 3AND

* plots
.plot v(Q) V(A) V(B) V(C)

* analasys
.tran 1n 60n




* main circuit file
.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 1

* * MUX test
Vdd Vdd 0 supplyVoltage

Va A 0 0
Vb B 0 0
Vc C 0 supplyVoltage

VS1 S1 0 PULSE(0, supplyVoltage, 13n, 1n, 1n, 7n, 20n)
VS2 S2 0 PULSE(0, supplyVoltage, 10n, 1n, 1n, 10n, 30n)

xMUX A B C S1 S2 OUT Vdd 0 MUX

* plots
.plot v(OUT) v(S1) v(S2)
.plot v(OUT)

* analasys
.tran 1n 60n




.param L = 0.1u
.param W = 10u

* NOT gate
.subckt NOT A Q Vdd Vss
   xMP1 Q A Vdd Vdd pmos1v l=L w=W
   xMN2 Q A Vss Vss nmos1v l=L w=W
.ends NOT

* NAND gate
.subckt NAND A B Q Vdd Vss
   * PMOS section
   xMP1 Vdd A Q Vdd pmos1v l=L w=W
   xMP2 Vdd B Q Vdd pmos1v l=L w=W

   * NMOS section
   xMN1 Q B 1 1 nmos1v l=L w=W
   xMN2 1 A Vss Vss nmos1v l=L w=W
.ends NAND

* AND gate
.subckt AND A B Q Vdd Vss
   xNAND A B intermediate Vdd Vss NAND
   xNOT intermediate Q Vdd Vss NOT
.ends



* main circuit file
.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 0.4

* MUX test
Vdd Vdd 0 supplyVoltage

Va A 0 0
Vb B 0 0
Vc C 0 supplyVoltage

V_D D 0 PULSE(0, supplyVoltage, 4n, 1n, 1n, 4n, 13n)
V_CLK CLK 0 PULSE(0, supplyVoltage, 0n, 1n, 1n, 10n, 20n)

xD_FLIP_FLOP D Q CLK Vdd 0 D_FLIP_FLOP

* plots
.plot v(Q) v(D) v(CLK)
.plot v(Q)
.plot v(CLK)
.plot v(D)

* analasys
.tran 1n 60n
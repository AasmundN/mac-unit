* MUX subcircuit
.subckt MUX A B S OUT Vdd Vss
   xAND1 S A 2 Vdd Vss AND
   xAND2 1 B 3 Vdd Vss AND

   xOR 2 3 OUT Vdd Vss OR

   xNOT S 1 Vdd Vss NOT
.ends
[aimspice]
[description]
448
* main circuit file
*.option gmin=1e-39

* includes
.include includes.cir

* params
.param supplyVoltage = 1
.param GND = 0

* circuit
Vdd Vdd GND supplyVoltage
R1 OUT GND 1k
V_CONTROL CONTROL GND PULSE(0, supplyVoltage, 0, 1n, 1n, 20n, 40n)
V_IN IN GND PULSE(0, supplyVoltage, 10n, 1n, 1n, 10n, 20n)

xTRANSMISSIONGATE IN OUT CONTROL Vdd GND TRANSMISSIONGATE

* plots
.plot V(IN) V(OUT) V(CONTROL)  

* analasys
*.tran 1n 60n
[tran]
1
60
X
X
0
[ana]
4 0
[end]

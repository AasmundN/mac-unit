* MUX subcircuit
.subckt MUX A B S OUT Vdd Vss
   * transmission gates
   xTRANSMISSION_GATEIN1 A OUT S NOT_S Vdd Vss TRANSMISSION_GATE 
   xTRANSMISSION_GATEIN2 B OUT NOT_S S Vdd Vss TRANSMISSION_GATE 

   * create inverted S
   xNOT S NOT_S Vdd Vss NOT
.ends
module multiplier(input bit a, input bit b, output bit out);
    assign out = a & b;
endmodule
